* C:\Users\lenovo\OneDrive\Desktop\project\q2.sch

* Schematics Version 9.1 - Web Update 1
* Thu Jun 16 18:08:18 2022



** Analysis setup **
.tran 7ms 10 0 2ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "q2.net"
.INC "q2.als"


.probe


.END
